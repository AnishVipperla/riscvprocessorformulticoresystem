module imm_decode (
    ports
);
    
endmodule