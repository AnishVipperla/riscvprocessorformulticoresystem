module alu (
    ports
);
    
endmodule